module Dec7s(a,q);
input [3:0] a;
output [7:0] q;
reg [7:0] q;
always @(a)
	begin 
	case(a)
		0:q=8'b11000000; 1:q=8'b11111001;
		2:q=8'b10100100; 3:q=8'b10110000;
		4:q=8'b10011001; 5:q=8'b10010010;
		6:q=8'b10000010; 7:q=8'b11111000;
		8:q=8'b10000000; 9:q=8'b10010000;
		10:q=8'b10001000; 11:q=8'b01111100;
		12:q=8'b00111001; 13:q=8'b01011110;
		14:q=8'b01111001; 15:q=8'b01110001;
	endcase
   end
endmodule 